module TOP(
    input A,
    input B,
    output F
);
    top U(.a(A),.b(B),.f(F) );
endmodule